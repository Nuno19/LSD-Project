library verilog;
use verilog.vl_types.all;
entity Proj_demo_vlg_vec_tst is
end Proj_demo_vlg_vec_tst;
